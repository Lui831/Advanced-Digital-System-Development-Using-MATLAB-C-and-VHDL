
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity Counter_syc is
    port (
        clk     : in  std_logic;
        reset   : in  std_logic;
        enable  : in  std_logic;
        count   : out std_logic_vector(3 downto 0)
    );
end entity Counter_syc;     



architecture Behavioral of Counter_syc is
    signal counter_reg : unsigned(3 downto 0) := (others => '0');   


process_counter:  process(clk, reset)
    begin       
        if clk'event and clk = '1' then
           if reset = '1' then
                counter_reg <= (others => '0');   
            elsif enable = '1' then
                counter_reg <= counter_reg + 1;   
            end if;
        end if;
    end process process_counter;    

  count <= std_logic_vector(counter_reg);     